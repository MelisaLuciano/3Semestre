��  CCircuit��  CSerializeHack           ��  CPart              ���  CEarth�� 	 CTerminal  � �      '           ��!f��=?    ��         ��      �� 	 CResistor��  CValue  k� ��     2k          @�@      �?k  
�  �� ��       +   ��#�?��!f��=?  
�  �� ��      '           ��!f��=�    �� ��          ��      ��  � 0�     1k        @�@      �?k  
�  ,� A�      +   ��#�?E\F5��M�  
�   � �      ,   ���^��?E\F5��M?    � ,�         ��      ��  CSPST��  CToggle  Pp8        
�  H4II     (    ��6k.?�k��=�  
�  HI      $    ��6k.?�k��=?    DL4         ��    ��  #� C�     2k          @�@      �?k  
�  H� I�       +   ��#�?�k��=?  
�  H� I�      $    ��6k.?�k��=�    D� L�          ��      ��    8          
�  �4�I     (    ��6k.?          
�  ��      %   ���^��?            ��4    "      ��    ��  �� ��     2k          @�@      �?k  
�  �� ��       ,   ���^��?          
�  �� ��      %   ���^��?            �� ��      &    ��      ��  �� ��     1k        @�@      �?k  
�  �� ��      ,   ���^��?@\F5��M�  
�  �� ��      -   Ǔ��@@\F5��M?    �� ��     *    ��      ��  �� ��     2k          @�@      �?k  
�  �� ��       -   Ǔ��@�2WV?  
�  �� ��      &    ��6k.?�2WV�    �� ��      .    ��      ��  ��8     0   
�  �4�I     (    ��6k.?�2WV�  
�  ��      &    ��6k.?�2WV?    ��4    2     ��    ��  p� ��     1k        @�@      �?k  
�  �� ��      -   Ǔ��@��0��b�  
�  `� u�      #         @��0��b?    t� ��     6    ��      ��  CBattery�  �)7    5V(          @      �? V 
�  ()%      #         @��Sk[�s�  
�  (<)Q     "           ��Sk[�s?    $4<     ;    ��      �
�  (`)u      "           ��Sk[�s�    t3|     >    ��      �� 
 CVoltmeter��  CMeter  ���    -4.32(    
�   x!�      *  ��?RE�          
�   �!�                             �,�     C    ��      �
�   �!�                              �+�     F    ��      ��  C741��  COpampSupply�� 
 CDummyPart  ����    K�  ����      ����    9V            "@      �? V       "�      �? V H 
�  ����     (    ��6k.?          
�  ����     !                     
�  ����     *  ��?RE����$��q?    ����     N      ��    �
�  ����      !                       ����     R    ��      ��  �^�l    1k        @�@      �?k  
�  �p�q     *  ��?RE�!��$��q�  
�  �p�q     (    ��6k.?!��$��q?    �l�t    U    ��      ��  3� S�     2k          @�@      �?k  
�  X� Y�       #         @N@w��zd?  
�  X� Y�      )    ��6k.?N@w��zd�    T� \�      Y    ��      ��  `�8     [   
�  X4YI     (    ��6k.?N@w��zd�  
�  XY      )    ��6k.?N@w��zd?    T\4    ]     ��    ?�A�  S�{�    -1.10(    
�  ����        B�����          
�  ����                            |���     a    ��      �
�  ����                             {���     d    ��      ��  n8|    1004        `�@      �?   
�  4�I�       B�����c�2��Q�  
�  ��        �t���?�c�2��Q?    |4�    g    ��      G�I�K�   �@�    K�   �@�      ��    9V            "@      �? V       "�      �? V i 
�  ��        �t���?          
�  ��                          
�  4�I�       B�������2��Q?    �4�     m      ��    �
�   ��                             � ��     q    ��      �
�  � h� }                 �c�2��Q�    � |� �     s    ��      ��  �� ��     32k          @�@      �?k  
�  �� ��       	   ffffff
@          
�  �� �	        ffffff
@            �� ��      v    ��      ��  �� �     64k          @�@      �?k  
�  � 	�       	   ffffff
@�#�Fz?  
�  � 		        �t���?�#�Fz�    � �      z    ��      ��  � ;�     128k          @�@      �?k  
�  @� A�       	   ffffff
@          
�  @� A	        ffffff
@            <� D�      ~    ��      ��  S� s�     256k          @A      �?k  
�  x� y�       	   ffffff
@�#�Fz�>  
�  x� y	        �t���?�#�Fz�    t� |�      �    ��      ��  s� ��     16k          @�@      �?k  
�  �� ��       	   ffffff
@�#�Fz+?  
�  �� �	        �t���?�#�Fz+�    �� ��      �    ��      ��  ;� [�     8k          @�@      �?k  
�  `� a�       	   ffffff
@          
�  `� a	        ffffff
@            \� d�      �    ��      ��  � #�     4k          @�@      �?k  
�  (� )�       	   ffffff
@�#�FzK?  
�  (� )	        �t���?�#�FzK�    $� ,�      �    ��      ��  � � � �     2k          @�@      �?k  
�  � � � �       	   ffffff
@          
�  � � � 	     
   ffffff
@            � � � �      �    ��      8��  k 1� ?    3.3V(    ffffff
@      �? V 
�  � � -      	   ffffff
@�c�2��Q�  
�  � D� Y                �c�2��Q?    � ,� D     �    ��      ��  (0H     �   
�  D	Y        �t���?�#�Fz�  
�  	-         �t���?�#�Fz?    ,D    �     ��    ��  �(�H      �   
�  �D�Y        �t���?          
�  ��-         ffffff
@            �,�D    �      ��    ��  H(hH      �   
�  @DAY        �t���?          
�  @A-         ffffff
@            <,DD    �      ��    ��  �(�H     �   
�  xDyY        �t���?�#�Fz�  
�  xy-         �t���?�#�Fz�>    t,|D    �     ��    ��  �(�H     �   
�  �D�Y        �t���?�#�Fz+�  
�  ��-         �t���?�#�Fz+?    �,�D    �     ��    ��  h(�H      �   
�  `DaY        �t���?          
�  `a-         ffffff
@            \,dD    �      ��    ��  � (H      �   
�  � D� Y        �t���?          
�  � � -      
   ffffff
@            � ,� D    �      ��    ��  0(PH     �   
�  (D)Y        �t���?�#�FzK�  
�  ()-         �t���?�#�FzK?    $,,D    �     ��                  ���  CWire  �� �      ' ��  ����     ( ��  x���     ( ��  xHy�      ( ��  XHyI     ( ��  xH�I     ( ��  �HII     ( ��  �H�I     ( ��  (� Y�      # ��  (� )      # ��  H� ��      + ��  @� I�      + ��  �� �      , ��  H� I	      $ ��  �� ��      , ��  �� ��      - ��  �� �	      % ��  �� ��      - ��  X� a�      # ��  �� �	      & ��  (P)a      " ��   p!y      * ��  �p!q     * ��   �!�        ��  ����     * ��  ����     ! ��  ����      ! ��  �p��      ( ��  �p�q     ( ��  �p�q     * ��  �p��      * ��  X� Y	      ) ��  ����       ��  P���      ��  ����       ��  � �� �       ��  � �� �      ��  � X� �       ��  H�Q�      ��  H�Q�      ��  � �	�      ��   �	�      ��   ��       ��  P�Q�       ��  � �	�      ��  (XaY      ��  � X� i       ��  �X�Y      ��  `X�Y      ��  @XyY      ��  XAY      ��  �X	Y      ��  � X)Y      ��  ��       ��  xy       ��  @A       ��  	       ��  ��       ��  `a       ��  ()       ��  � �       
 ��  @� y�      	 ��  � A�      	 ��  �� 	�      	 ��  �� ��      	 ��  `� ��      	 ��  (� a�      	 ��  � � )�      	 ��  � � � �      	 ��  � � �       	               �                             �   �    �   �  �    �  �   �    � " " � # � # & � & ' ' � * * � + � + . � . / / � 2 2 � 3 � 3 6 6 � 7 � 7 ; � ; < < � > � > C � C D D � F � F J J N � N O � O P P � R � R U U � V � V Y � Y Z Z � ] ] � ^ � ^ a � a b b � d � d g g � h � h j j m � m n � n o o � q � q s � s v � v w w � z � z { { � ~ � ~   � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �   � N � � � � ] � � � "  2 � � Y � ; �    &    * � . + ' # 6 � � 7 / 3 < > � C � � D F P � � O � R � � � V U � � � Z ^ � a � � b d � � � � � � o � g � � h � n � q � � � m � � � s � � � � � � � � � � � � � � � �  � { � w � � � � � � � ~ � z � � � � v � � � � � � � � � �  .          �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 